jesper@dhcp-073151.eduroam.chalmers.se.947